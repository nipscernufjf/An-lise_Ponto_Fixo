library verilog;
use verilog.vl_types.all;
entity procm6_tb is
end procm6_tb;
